module ASIP()
endmodule
