module ASIP()

