module Vector_Mux_8 #(I=20,L=8)(input  [3:0]   			S,
										  input  [I-1:0][L-1:0] D08, D09, D10, D11, D12, D13, D14, D15,
										  output [I-1:0][L-1:0] Y);

logic[I-1:0][L-1:0] out;	
							
always_comb begin
	case(S)
		4'b1000: out = D08;
		4'b1001: out = D09;
		4'b1010: out = D10; 
		4'b1011: out = D11;
		4'b1100: out = D12;
		4'b1101: out = D13;
		4'b1110: out = D14;
		4'b1111: out = D15;
		default: out = 0;
	endcase
end

assign Y = out;

endmodule