module ASIP();

endmodule