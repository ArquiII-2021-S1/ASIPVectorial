module ASIP();
    
endmodule
